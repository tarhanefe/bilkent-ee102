library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
----------------------------
-- 0 => BEGIN
-- 1 => END
----------------------------
entity GAME_END_BEGIN_W is
PORT(
SEL_END_BEGIN : in STD_LOGIC;
CLR : in STD_LOGIC;
VIDON: in STD_LOGIC;
HC : in STD_LOGIC_VECTOR(10 downto 0);
VC : in STD_LOGIC_VECTOR(10 downto 0);
RED : out STD_LOGIC_VECTOR(3 downto 0);
GREEN : out STD_LOGIC_VECTOR(3 downto 0);
BLUE : out STD_LOGIC_VECTOR(3 downto 0)
);
end GAME_END_BEGIN_W;

architecture GAME_END_BEGIN_W of GAME_END_BEGIN_W is
SIGNAL R : STD_LOGIC_VECTOR(71 DOWNTO 0); 
SIGNAL G : STD_LOGIC_VECTOR(71 DOWNTO 0); 
SIGNAL B : STD_LOGIC_VECTOR(71 DOWNTO 0); 
SIGNAL R1,R2,R3,R4,R5,R6,R7,R8,R9,R10,R11 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL B1,B2,B3,B4,B5,B6,B7,B8,B9,B10,B11 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11 : STD_LOGIC_VECTOR(3 DOWNTO 0);
CONSTANT A : INTEGER := 10;
COMPONENT WORD_SELECTOR
PORT(
SEL_WORD : in std_logic_vector(7 downto 0);
R : in integer:= 0;
C : in integer:= 0;
HC : in STD_LOGIC_VECTOR (10 downto 0);
VC : in STD_LOGIC_VECTOR (10 downto 0);
RED : out STD_LOGIC_VECTOR (3 downto 0);
GREEN : out STD_LOGIC_VECTOR (3 downto 0);
BLUE : out STD_LOGIC_VECTOR (3 downto 0)
);

END COMPONENT;

COMPONENT CHAR_PLACER
PORT(
MUX_IN: in STD_LOGIC_VECTOR(7 downto 0);
R : in integer;
C : in integer;
HC : in STD_LOGIC_VECTOR (10 downto 0);
VC : in STD_LOGIC_VECTOR (10 downto 0);
RED : out STD_LOGIC_VECTOR (3 downto 0);
GREEN : out STD_LOGIC_VECTOR (3 downto 0);
BLUE : out STD_LOGIC_VECTOR (3 downto 0));
END COMPONENT;
begin
---------------------------------------------

UM1: CHAR_PLACER
PORT MAP(
MUX_IN => x"16",
R => 120,
C => 224-A,
HC => HC,
VC => VC,
RED => R1,
GREEN => G1,
BLUE => B1
);
UM2: CHAR_PLACER
PORT MAP(
MUX_IN => x"07",
R => 120,
C => 232-A,
HC => HC,
VC => VC,
RED => R2,
GREEN => G2,
BLUE => B2
);
UM3: CHAR_PLACER
PORT MAP(
MUX_IN => x"00",
R => 120,
C => 240-A,
HC => HC,
VC => VC,
RED => R3,
GREEN => G3,
BLUE => B3
);
UM4: CHAR_PLACER
PORT MAP(
MUX_IN => x"02",
R => 120,
C => 248-A,
HC => HC,
VC => VC,
RED => R4,
GREEN => G4,
BLUE => B4
);
UM5: CHAR_PLACER
PORT MAP(
MUX_IN => x"0A",
R => 120,
C => 256-A,
HC => HC,
VC => VC,
RED => R5,
GREEN => G5,
BLUE => B5
);
UM6: CHAR_PLACER
PORT MAP(
MUX_IN => x"25",
R => 120,
C => 264-A,
HC => HC,
VC => VC,
RED => R6,
GREEN => G6,
BLUE => B6
);
UM7: CHAR_PLACER
PORT MAP(
MUX_IN => x"00",
R => 120,
C => 272-A,
HC => HC,
VC => VC,
RED => R7,
GREEN => G7,
BLUE => B7
);

UM8: CHAR_PLACER
PORT MAP(
MUX_IN => x"25",
R => 120,
C => 280-A,
HC => HC,
VC => VC,
RED => R8,
GREEN => G8,
BLUE => B8
);
UM9: CHAR_PLACER
PORT MAP(
MUX_IN => x"0C",
R => 120,
C => 288-A,
HC => HC,
VC => VC,
RED => R9,
GREEN => G9,
BLUE => B9
);
UM10: CHAR_PLACER
PORT MAP(
MUX_IN => x"0E",
R => 120,
C => 296-A,
HC => HC,
VC => VC,
RED => R10,
GREEN => G10,
BLUE => B10
);

UM11: CHAR_PLACER
PORT MAP(
MUX_IN => x"0B",
R => 120,
C => 304-A,
HC => HC,
VC => VC,
RED => R11,
GREEN => G11,
BLUE => B11
);
U1: CHAR_PLACER
PORT MAP(
MUX_IN => x"04",
R => 120,
C => 312-A,
HC => HC,
VC => VC,
RED => R(71 DOWNTO 68),
GREEN => G(71 DOWNTO 68),
BLUE => B(71 DOWNTO 68)
);
----------------------------------------------
U2: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"07",
R => 120,
C => 328-A,
HC => HC,
VC => VC,
RED => R(67 DOWNTO 64),
GREEN => G(67 DOWNTO 64),
BLUE => B(67 DOWNTO 64)
);

U3: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"0C",
R => 120,
C => 368-A,
HC => HC,
VC => VC,
RED => R(63 DOWNTO 60),
GREEN => G(63 DOWNTO 60),
BLUE => B(63 DOWNTO 60)
);

U4: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"0A",
R => 120,
C => 392-A,
HC => HC,
VC => VC,
RED => R(59 DOWNTO 56),
GREEN => G(59 DOWNTO 56),
BLUE => B(59 DOWNTO 56)
);

U5: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"03",
R => 120,
C => 424-A,
HC => HC,
VC => VC,
RED => R(55 DOWNTO 52),
GREEN => G(55 DOWNTO 52),
BLUE => B(55 DOWNTO 52)
);
-------------------------------------------------------
U6: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"05",
R => 360,
C => 240,
HC => HC,
VC => VC,
RED => R(51 DOWNTO 48),
GREEN => G(51 DOWNTO 48),
BLUE => B(51 DOWNTO 48)
);

U7: CHAR_PLACER
PORT MAP(
MUX_IN => x"28",
R => 360,
C => 288,
HC => HC,
VC => VC,
RED => R(47 DOWNTO 44),
GREEN => G(47 DOWNTO 44),
BLUE => B(47 DOWNTO 44)
);

U8: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"0B",
R => 360,
C => 304,
HC => HC,
VC => VC,
RED => R(43 DOWNTO 40),
GREEN => G(43 DOWNTO 40),
BLUE => B(43 DOWNTO 40)
);

U9: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"07",
R => 360,
C => 336,
HC => HC,
VC => VC,
RED => R(39 DOWNTO 36),
GREEN => G(39 DOWNTO 36),
BLUE => B(39 DOWNTO 36)
);

-----------------------------------------------------
U14: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"07",
R => 240,
C => 288,
HC => HC,
VC => VC,
RED => R(19 DOWNTO 16),
GREEN => G(19 DOWNTO 16),
BLUE => B(19 DOWNTO 16)
);

U15: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"12",
R => 240,
C => 328,
HC => HC,
VC => VC,
RED => R(15 DOWNTO 12),
GREEN => G(15 DOWNTO 12),
BLUE => B(15 DOWNTO 12)
);
--------------------------------
U16: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"04",
R => 360,
C => 256,
HC => HC,
VC => VC,
RED => R(11 DOWNTO 8),
GREEN => G(11 DOWNTO 8),
BLUE => B(11 DOWNTO 8)
);

U17: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"0B",
R => 360,
C => 312,
HC => HC,
VC => VC,
RED => R(7 DOWNTO 4),
GREEN => G(7 DOWNTO 4),
BLUE => B(7 DOWNTO 4)
);

U18: WORD_SELECTOR
PORT MAP(
SEL_WORD => x"01",
R => 360,
C => 344,
HC => HC,
VC => VC,
RED => R(3 DOWNTO 0),
GREEN => G(3 DOWNTO 0),
BLUE => B(3 DOWNTO 0)
);
-------------------------------------
PROCESS(VIDON,SEL_END_BEGIN,R,G,B)
BEGIN
CASE SEL_END_BEGIN IS
WHEN '0' => --- BEGIN SCREEN
IF VIDON = '1' THEN
RED <= R(71 DOWNTO 68) OR R(67 DOWNTO 64) OR R(63 DOWNTO 60) OR R(59 DOWNTO 56) OR R(55 DOWNTO 52) OR R(51 DOWNTO 48) OR R(47 DOWNTO 44) OR R(43 DOWNTO 40) OR R(39 DOWNTO 36)
OR R1 OR R2 OR R3 OR R4 OR R5 OR R6 OR R7 OR R8 OR R9 OR R10 OR R11;
GREEN <= X"0" OR G(67 DOWNTO 64) OR G(63 DOWNTO 60) OR G(59 DOWNTO 56) OR G(55 DOWNTO 52) OR G(51 DOWNTO 48) OR G(47 DOWNTO 44) OR G(43 DOWNTO 40) OR G(39 DOWNTO 36)
OR G1 OR G2 OR G3 OR G4 OR G5 OR G6 OR G7 OR G8 OR X"0" OR X"0" OR X"0";
BLUE <= B(71 DOWNTO 68) OR B(67 DOWNTO 64) OR B(63 DOWNTO 60) OR B(59 DOWNTO 56) OR B(55 DOWNTO 52) OR B(51 DOWNTO 48) OR B(47 DOWNTO 44) OR B(43 DOWNTO 40) OR B(39 DOWNTO 36)
OR X"0" OR X"0" OR X"0" OR X"0" OR X"0" OR B6 OR B7 OR B8 OR B9 OR B10 OR B11;
ELSE 
RED <= "0000";
GREEN <= "0000";
BLUE <= "0000";
END IF;

WHEN '1' =>  ----ENDING SCREEN
IF VIDON = '1' THEN
RED <= R(19 DOWNTO 16) OR R(15 DOWNTO 12) OR R(11 DOWNTO 8) OR R(7 DOWNTO 4) OR R(3 DOWNTO 0);
GREEN <= G(19 DOWNTO 16) OR G(15 DOWNTO 12) OR G(11 DOWNTO 8) OR G(7 DOWNTO 4) OR G(3 DOWNTO 0);
BLUE <= B(19 DOWNTO 16) OR B(15 DOWNTO 12) OR B(11 DOWNTO 8) OR B(7 DOWNTO 4) OR B(3 DOWNTO 0);
ELSE 
RED <= "0000";
GREEN <= "0000";
BLUE <= "0000";
END IF;

END CASE;
END PROCESS;


end GAME_END_BEGIN_W;