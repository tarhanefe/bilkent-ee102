library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
--------------------------------
entity SCORE_COUNT is
PORT(
DIF : IN STD_LOGIC;
CLK : IN STD_LOGIC;
RESET : IN STD_LOGIC;
BTN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
GAME_OVER : OUT STD_LOGIC;
SQUARES : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
SCORE : OUT INTEGER:= 0
);
end SCORE_COUNT;
--------------------------------
architecture Behavioral of SCORE_COUNT is
TYPE STATE_TYPE IS (S_CATCH,S_MISS,S_OVER,S_INIT,S_WAIT);
SIGNAL MOLE : STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL STATE : STATE_TYPE;
SIGNAL SCOREE : INTEGER := 5;
SIGNAL RAND : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL BTN0P,BTN0R,BTN1P,BTN1R,BTN2P,BTN2R,BTN3P,BTN3R,BTN4P,BTN4R : STD_LOGIC;
SIGNAL CLK_G,CLK_W : STD_LOGIC;
SIGNAL PUSHED : STD_LOGIC;
------------------------------------
COMPONENT LFSR4 IS
PORT(
DIF : IN STD_LOGIC;
CLK : IN STD_LOGIC;
RAND_COLOR : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
RAND_NUMB : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
END COMPONENT;
-----------------------
COMPONENT PUSH_RELEASE IS
PORT(
CLK : IN STD_LOGIC;
BTN_IN : IN STD_LOGIC;
BTN_OUT_P : OUT STD_LOGIC;
BTN_OUT_R : OUT STD_LOGIC
);
END COMPONENT;

---------------------------
BEGIN
RANDOM_GEN : LFSR4 
PORT MAP(
DIF => DIF,
CLK => CLK,
RAND_COLOR => MOLE,
RAND_NUMB => RAND
);
------------------------------
BTN0 : PUSH_RELEASE PORT MAP(CLK => CLK, BTN_IN => BTN(0),BTN_OUT_P => BTN0P,BTN_OUT_R => BTN0R );
BTN1 : PUSH_RELEASE PORT MAP(CLK => CLK, BTN_IN => BTN(1),BTN_OUT_P => BTN1P,BTN_OUT_R => BTN1R );
BTN2 : PUSH_RELEASE PORT MAP(CLK => CLK, BTN_IN => BTN(2),BTN_OUT_P => BTN2P,BTN_OUT_R => BTN2R );
BTN3 : PUSH_RELEASE PORT MAP(CLK => CLK, BTN_IN => BTN(3),BTN_OUT_P => BTN3P,BTN_OUT_R => BTN3R );
BTN4 : PUSH_RELEASE PORT MAP(CLK => CLK, BTN_IN => BTN(4),BTN_OUT_P => BTN4P,BTN_OUT_R => BTN4R );
PUSHED <= BTN0P OR BTN1P OR BTN2P OR BTN3P OR BTN4P;
SQUARES <= MOLE;
SCORE <= SCOREE;
-----------------------
PROCESS(CLK)
VARIABLE CAUGHT : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
IF RESET = '1' THEN
STATE <= S_INIT;
ELSIF RISING_EDGE(CLK) THEN
CASE STATE IS

WHEN S_INIT =>
GAME_OVER <= '0';
SCOREE <= 10;
IF BTN0P = '1' THEN
STATE <= S_WAIT;
ELSE
STATE <= S_INIT;
END IF;
------------------------------------
WHEN S_WAIT =>
IF SCOREE > 0 THEN
IF PUSHED /= '0' THEN
IF BTN = MOLE AND CAUGHT /= RAND THEN
STATE <= S_CATCH;
ELSIF BTN /= MOLE THEN
STATE <= S_MISS; 
END IF;
ELSE
STATE <= S_WAIT;
END IF;
ELSE
STATE <= S_OVER;
END IF;
------------------------------------
WHEN S_MISS => 
SCOREE <= SCOREE - 1;
CAUGHT := RAND;
STATE <= S_WAIT;
------------------------------------
WHEN S_CATCH => 
SCOREE <= SCOREE + 1;
CAUGHT := RAND;
STATE <= S_WAIT;
------------------------------------
WHEN S_OVER =>
GAME_OVER <= '1';
STATE <= S_OVER;
------------------------------------
END CASE;
END IF;
END PROCESS;
end Behavioral;
