library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
------------------------------
ENTITY RANDOM_CLK_DIV is
PORT (  
DIF : IN STD_LOGIC;
CLK : in std_logic;
CLK_O : out std_logic);		  
end RANDOM_CLK_DIV;
-----------------------------
ARCHITECTURE RANDOM_CLK_DIV of RANDOM_CLK_DIV is
CONSTANT COUNT1 : INTEGER := (17500000);  
CONSTANT COUNT2 : INTEGER := (25000000);
SIGNAL COUNT : INTEGER := (17500000);
SIGNAL TMP : std_logic := '0'; 
------------------------------
BEGIN
PROCESS(CLK,DIF)
BEGIN 
IF RISING_EDGE(CLK) THEN
CASE DIF IS
WHEN '0' => COUNT <= COUNT1;
WHEN '1' => COUNT <= COUNT2;
END CASE;
END IF;
END PROCESS;
DIV_CLK: PROCESS(CLK,TMP)              
VARIABLE DIV_CNT : integer := 0;   
BEGIN
IF (rising_edge(clk)) THEN   
IF (DIV_CNT = COUNT) THEN
TMP <= NOT TMP; 
DIV_CNT := 0; 
ELSIF DIV_CNT < COUNT THEN
DIV_CNT := DIV_CNT + 1; 
ELSE
DIV_CNT := 0;
END IF; 
END IF; 
CLK_O <= TMP; 
END PROCESS DIV_CLK; 
END RANDOM_CLK_DIV;